package apb_pkg;                       // package declaration
  
  import uvm_pkg::*; 
  `include "uvm_macros.svh"                  // import UVM package
`include "sequence_item.sv"
`include "seque.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "env.sv"
`include "apb_test.sv"
  
endpackage 
